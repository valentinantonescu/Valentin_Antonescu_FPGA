module transcodor (input [4:0] s,
						 output reg [13:0] q);
	
			always@(s)
				case(s)
					  5'b00000: q=14'b10000001000000; //0
				     5'b00001: q=14'b10000001111001; //1
					  5'b00010: q=14'b10000000100100; //2
					  5'b00011: q=14'b10000000110000; //3
					  5'b00100: q=14'b10000001111001; //4
					  5'b00101: q=14'b10000000010010; //5
					  5'b00110: q=14'b10000000000010; //6
					  5'b00111: q=14'b10000001111000; //7
					  5'b01000: q=14'b10000000100100; //8
					  5'b01001: q=14'b10000000010000; //9
					  5'b01010: q=14'b11110011000000; //10
					  5'b01011: q=14'b11110011111001; //11
					  5'b01100: q=14'b10000000110000; //12
					  5'b01101: q=14'b11110010110000; //13
					  5'b01110: q=14'b11110010011001; //14
					  5'b01111: q=14'b11110010010010; //15
					  5'b10000: q=14'b10000000011001; //16
				     5'b10001: q=14'b11110011111000; //17
					  5'b10010: q=14'b11110010000000; //18
					  5'b10011: q=14'b11110010010000; //19
					  5'b10100: q=14'b10000000010010; //20
					  5'b10101: q=14'b01001001111001; //21
					  5'b10110: q=14'b01001000100100; //22
					  5'b10111: q=14'b01001000110000; //23
					  5'b11000: q=14'b10000000000010; //24
					  5'b11001: q=14'b01001000010010; //25
					  5'b11010: q=14'b01001000000010; //26
					  5'b11011: q=14'b01001001111000; //27
					  5'b11100: q=14'b10000001111000; //28
					  5'b11101: q=14'b01001000010000; //29
					  5'b11110: q=14'b01100001000000; //30
					  5'b11111: q=14'b01100001111001; //31
					  default:  q=14'b10000001000000;
					  
				endcase
			
endmodule