module transcodor (input [6:0] s,
						 output reg [13:0] q);
	
			always@(s)
				case(s)
					  7'b0000000: q=14'b10000001000000; //0
					  7'b0000100: q=14'b10000001111001; //1
					  7'b0001000: q=14'b10000000100100; //2
					  7'b0001100: q=14'b10000000110000; //3
					  7'b0010000: q=14'b10000000011001; //4
					  7'b0010100: q=14'b10000000010010; //5
					  7'b0011000: q=14'b10000000000010; //6
					  7'b0011100: q=14'b10000001111000; //7
					  7'b0100000: q=14'b10000000000000; //8
					  7'b0100100: q=14'b10000000010000; //9
					  7'b0101000: q=14'b11110011000000; //10
					  7'b0101100: q=14'b11110011111001; //11
					  7'b0110000: q=14'b11110010100100; //12
					  7'b0110100: q=14'b11110010110000; //13
					  7'b0111000: q=14'b11110010011001; //14
					  7'b0111100: q=14'b11110010010010; //15
					  7'b1000000: q=14'b11110010000010; //16
					  7'b1000100: q=14'b11110011111000; //17
					  7'b1001000: q=14'b11110010000000; //18
					  7'b1001100: q=14'b11110010010000; //19
					  7'b1010000: q=14'b01001001000000; //20
					  7'b1010100: q=14'b01001001111001; //21
					  7'b1011000: q=14'b01001000100100; //22
					  7'b1011100: q=14'b01001000110000; //23
					  7'b1100000: q=14'b01001000011001; //24
					  7'b1100100: q=14'b01001000010010; //25
					  7'b1101000: q=14'b01001000000010; //26
					  7'b1101100: q=14'b01001001111000; //27
					  7'b1110000: q=14'b01001000000000; //28
					  7'b1110100: q=14'b01001000010000; //29
					  7'b1111000: q=14'b01100001000000; //30
					  7'b1111100: q=14'b01100001111001; //31
					  default:    q=14'b10000001111001;
					  
				endcase
			
endmodule