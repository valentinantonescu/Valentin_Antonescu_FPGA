module slave_I2C