module transcodor (input [3:0] s,
						 output reg [6:0] q);
	
			always@(s)
				case(s)
					  4'b0000: q=7'b1000000;
				          4'b0001: q=7'b1111001;
					  4'b0010: q=7'b0100100;
					  4'b0011: q=7'b0110000;
					  4'b0100: q=7'b0011001;
					  4'b0101: q=7'b0010010;
					  4'b0110: q=7'b0000010;
					  4'b0111: q=7'b1111000;
					  4'b1000: q=7'b0000000;
					  4'b1001: q=7'b0010000;
					  4'b1010: q=7'b0001000;
					  4'b1011: q=7'b0000011;
					  4'b1100: q=7'b1000110;
					  4'b1101: q=7'b0100001;
					  4'b1110: q=7'b0000110;
					  4'b1111: q=7'b0001110;
					  
				endcase
			
endmodule
