module master_I2C